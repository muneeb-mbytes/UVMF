//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
// This file contains defines and typedefs to be compiled for use in
// the simulation running on the host server when using Veloce.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
`ifndef TYPEDEFS_HVL
`definr TYPEDEFS_HVL

// pragma uvmf custom additional begin
// pragma uvmf custom additional end
`endif
