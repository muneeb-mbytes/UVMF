//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: This class defines the variables required for an wishbone_slave
//    transaction.  Class variables to be displayed in waveform transaction
//    viewing are added to the transaction viewing stream in the add_to_wave
//    function.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
class wishbone_slave_transaction  extends uvmf_transaction_base;

  `uvm_object_utils( wishbone_slave_transaction )

  bit sck ;
  rand bit cs ;
  rand bit mosi ;
  bit miso ;

  //Constraints for the transaction variables:

  // pragma uvmf custom class_item_additional begin
  // pragma uvmf custom class_item_additional end

  //*******************************************************************
  //*******************************************************************
  // Macros that define structs and associated functions are
  // located in wishbone_slave_macros.svh

  //*******************************************************************
  // Monitor macro used by wishbone_slave_monitor and wishbone_slave_monitor_bfm
  // This struct is defined in wishbone_slave_macros.svh
  `wishbone_slave_MONITOR_STRUCT
    wishbone_slave_monitor_s wishbone_slave_monitor_struct;
  //*******************************************************************
  // FUNCTION: to_monitor_struct()
  // This function packs transaction variables into a wishbone_slave_monitor_s
  // structure.  The function returns the handle to the wishbone_slave_monitor_struct.
  // This function is defined in wishbone_slave_macros.svh
  `wishbone_slave_TO_MONITOR_STRUCT_FUNCTION 
  //*******************************************************************
  // FUNCTION: from_monitor_struct()
  // This function unpacks the struct provided as an argument into transaction 
  // variables of this class.
  // This function is defined in wishbone_slave_macros.svh
  `wishbone_slave_FROM_MONITOR_STRUCT_FUNCTION 

  //*******************************************************************
  // Initiator macro used by wishbone_slave_driver and wishbone_slave_driver_bfm
  // to communicate initiator driven data to wishbone_slave_driver_bfm.
  // This struct is defined in wishbone_slave_macros.svh
  `wishbone_slave_INITIATOR_STRUCT
    wishbone_slave_initiator_s wishbone_slave_initiator_struct;
  //*******************************************************************
  // FUNCTION: to_initiator_struct()
  // This function packs transaction variables into a wishbone_slave_initiator_s
  // structure.  The function returns the handle to the wishbone_slave_initiator_struct.
  // This function is defined in wishbone_slave_macros.svh
  `wishbone_slave_TO_INITIATOR_STRUCT_FUNCTION  
  //*******************************************************************
  // FUNCTION: from_initiator_struct()
  // This function unpacks the struct provided as an argument into transaction 
  // variables of this class.
  // This function is defined in wishbone_slave_macros.svh
  `wishbone_slave_FROM_INITIATOR_STRUCT_FUNCTION 

  //*******************************************************************
  // Responder macro used by wishbone_slave_driver and wishbone_slave_driver_bfm
  // to communicate Responder driven data to wishbone_slave_driver_bfm.
  // This struct is defined in wishbone_slave_macros.svh
  `wishbone_slave_RESPONDER_STRUCT
    wishbone_slave_responder_s wishbone_slave_responder_struct;
  //*******************************************************************
  // FUNCTION: to_responder_struct()
  // This function packs transaction variables into a wishbone_slave_responder_s
  // structure.  The function returns the handle to the wishbone_slave_responder_struct.
  // This function is defined in wishbone_slave_macros.svh
  `wishbone_slave_TO_RESPONDER_STRUCT_FUNCTION 
  //*******************************************************************
  // FUNCTION: from_responder_struct()
  // This function unpacks the struct provided as an argument into transaction 
  // variables of this class.
  // This function is defined in wishbone_slave_macros.svh
  `wishbone_slave_FROM_RESPONDER_STRUCT_FUNCTION 
  // ****************************************************************************
  // FUNCTION : new()
  // This function is the standard SystemVerilog constructor.
  //
  function new( string name = "" );
    super.new( name );
  endfunction

  // ****************************************************************************
  // FUNCTION: convert2string()
  // This function converts all variables in this class to a single string for 
  // logfile reporting.
  //
  virtual function string convert2string();
    // pragma uvmf custom convert2string begin
    // UVMF_CHANGE_ME : Customize format if desired.
    return $sformatf("sck:0x%x cs:0x%x mosi:0x%x miso:0x%x ",sck,cs,mosi,miso);
    // pragma uvmf custom convert2string end
  endfunction

  //*******************************************************************
  // FUNCTION: do_print()
  // This function is automatically called when the .print() function
  // is called on this class.
  //
  virtual function void do_print(uvm_printer printer);
    // pragma uvmf custom do_print begin
    // UVMF_CHANGE_ME : Current contents of do_print allows for the use of UVM 1.1d, 1.2 or P1800.2.
    // Update based on your own printing preference according to your preferred UVM version
    $display(convert2string());
    // pragma uvmf custom do_print end
  endfunction

  //*******************************************************************
  // FUNCTION: do_compare()
  // This function is automatically called when the .compare() function
  // is called on this class.
  //
  virtual function bit do_compare (uvm_object rhs, uvm_comparer comparer);
    wishbone_slave_transaction  RHS;
    if (!$cast(RHS,rhs)) return 0;
    // pragma uvmf custom do_compare begin
    // UVMF_CHANGE_ME : Eliminate comparison of variables not to be used for compare
    return (super.do_compare(rhs,comparer)
            &&(this.sck == RHS.sck)
            &&(this.cs == RHS.cs)
            &&(this.mosi == RHS.mosi)
            &&(this.miso == RHS.miso)
            );
    // pragma uvmf custom do_compare end
  endfunction

  //*******************************************************************
  // FUNCTION: do_copy()
  // This function is automatically called when the .copy() function
  // is called on this class.
  //
  virtual function void do_copy (uvm_object rhs);
    wishbone_slave_transaction  RHS;
    assert($cast(RHS,rhs));
    // pragma uvmf custom do_copy begin
    super.do_copy(rhs);
    this.sck = RHS.sck;
    this.cs = RHS.cs;
    this.mosi = RHS.mosi;
    this.miso = RHS.miso;
    // pragma uvmf custom do_copy end
  endfunction

  // ****************************************************************************
  // FUNCTION: add_to_wave()
  // This function is used to display variables in this class in the waveform 
  // viewer.  The start_time and end_time variables must be set before this 
  // function is called.  If the start_time and end_time variables are not set
  // the transaction will be hidden at 0ns on the waveform display.
  // 
  virtual function void add_to_wave(int transaction_viewing_stream_h);
    `ifdef QUESTA
    if (transaction_view_h == 0) begin
      transaction_view_h = $begin_transaction(transaction_viewing_stream_h,"wishbone_slave_transaction",start_time);
    end
    super.add_to_wave(transaction_view_h);
    // pragma uvmf custom add_to_wave begin
    // UVMF_CHANGE_ME : Color can be applied to transaction entries based on content, example below
    // case()
    //   1 : $add_color(transaction_view_h,"red");
    //   default : $add_color(transaction_view_h,"grey");
    // endcase
    // UVMF_CHANGE_ME : Eliminate transaction variables not wanted in transaction viewing in the waveform viewer
    $add_attribute(transaction_view_h,sck,"sck");
    $add_attribute(transaction_view_h,cs,"cs");
    $add_attribute(transaction_view_h,mosi,"mosi");
    $add_attribute(transaction_view_h,miso,"miso");
    // pragma uvmf custom add_to_wave end
    $end_transaction(transaction_view_h,end_time);
    $free_transaction(transaction_view_h);
    `endif // QUESTA
  endfunction

endclass

// pragma uvmf custom external begin
// pragma uvmf custom external end

