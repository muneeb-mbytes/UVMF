//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
// DESCRIPTION: Protocol specific agent class definition
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//

`ifndef SPI_S_AGENT
`define SPI_S_AGENT

class spi_s_agent  extends uvmf_parameterized_agent #(
                    .CONFIG_T(spi_s_configuration ),
                    .DRIVER_T(spi_s_driver ),
                    .MONITOR_T(spi_s_monitor ),
                    .COVERAGE_T(spi_s_transaction_coverage ),
                    .TRANS_T(spi_s_transaction )
                    );

  `uvm_component_utils( spi_s_agent )

// pragma uvmf custom class_item_additional begin
// pragma uvmf custom class_item_additional end

// ****************************************************************************
// FUNCTION : new()
// This function is the standard SystemVerilog constructor.
//
  function new( string name = "", uvm_component parent = null );
    super.new( name, parent );
  endfunction

// ****************************************************************************
  // FUNCTION: build_phase
  virtual function void build_phase(uvm_phase phase);
// pragma uvmf custom build_phase_pre_super begin
// pragma uvmf custom build_phase_pre_super end
    super.build_phase(phase);
    if (configuration.active_passive == ACTIVE) begin
      // Place sequencer handle into configuration object
      // so that it may be retrieved from configuration 
      // rather than using uvm_config_db
      configuration.sequencer = this.sequencer;
    end
  endfunction
  
endclass


// pragma uvmf custom external begin
// pragma uvmf custom external end
`endif
