//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: This class defines the variables required for an mem
//    transaction.  Class variables to be displayed in waveform transaction
//    viewing are added to the transaction viewing stream in the add_to_wave
//    function.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
class mem_transaction #(
      int DATA_WIDTH = 220,
      int ADDR_WIDTH = 210
      ) extends uvmf_transaction_base;

  `uvm_object_param_utils( mem_transaction #(
                           DATA_WIDTH,
                           ADDR_WIDTH
                           ))

  bit [DATA_WIDTH-1:0] read_data ;
  bit [DATA_WIDTH-1:0] write_data ;
  rand bit [ADDR_WIDTH-1:0] address ;
  rand bit [3:0] byte_enable ;
  int chksum ;

  //Constraints for the transaction variables:
  constraint address_word_align_c { address[1:0]==0; }

  // pragma uvmf custom class_item_additional begin
  // pragma uvmf custom class_item_additional end

  //*******************************************************************
  //*******************************************************************
  // Macros that define structs and associated functions are
  // located in mem_macros.svh

  //*******************************************************************
  // Monitor macro used by mem_monitor and mem_monitor_bfm
  // This struct is defined in mem_macros.svh
  `mem_MONITOR_STRUCT
    mem_monitor_s mem_monitor_struct;
  //*******************************************************************
  // FUNCTION: to_monitor_struct()
  // This function packs transaction variables into a mem_monitor_s
  // structure.  The function returns the handle to the mem_monitor_struct.
  // This function is defined in mem_macros.svh
  `mem_TO_MONITOR_STRUCT_FUNCTION 
  //*******************************************************************
  // FUNCTION: from_monitor_struct()
  // This function unpacks the struct provided as an argument into transaction 
  // variables of this class.
  // This function is defined in mem_macros.svh
  `mem_FROM_MONITOR_STRUCT_FUNCTION 

  //*******************************************************************
  // Initiator macro used by mem_driver and mem_driver_bfm
  // to communicate initiator driven data to mem_driver_bfm.
  // This struct is defined in mem_macros.svh
  `mem_INITIATOR_STRUCT
    mem_initiator_s mem_initiator_struct;
  //*******************************************************************
  // FUNCTION: to_initiator_struct()
  // This function packs transaction variables into a mem_initiator_s
  // structure.  The function returns the handle to the mem_initiator_struct.
  // This function is defined in mem_macros.svh
  `mem_TO_INITIATOR_STRUCT_FUNCTION  
  //*******************************************************************
  // FUNCTION: from_initiator_struct()
  // This function unpacks the struct provided as an argument into transaction 
  // variables of this class.
  // This function is defined in mem_macros.svh
  `mem_FROM_INITIATOR_STRUCT_FUNCTION 

  //*******************************************************************
  // Responder macro used by mem_driver and mem_driver_bfm
  // to communicate Responder driven data to mem_driver_bfm.
  // This struct is defined in mem_macros.svh
  `mem_RESPONDER_STRUCT
    mem_responder_s mem_responder_struct;
  //*******************************************************************
  // FUNCTION: to_responder_struct()
  // This function packs transaction variables into a mem_responder_s
  // structure.  The function returns the handle to the mem_responder_struct.
  // This function is defined in mem_macros.svh
  `mem_TO_RESPONDER_STRUCT_FUNCTION 
  //*******************************************************************
  // FUNCTION: from_responder_struct()
  // This function unpacks the struct provided as an argument into transaction 
  // variables of this class.
  // This function is defined in mem_macros.svh
  `mem_FROM_RESPONDER_STRUCT_FUNCTION 
  // ****************************************************************************
  // FUNCTION : new()
  // This function is the standard SystemVerilog constructor.
  //
  function new( string name = "" );
    super.new( name );
  endfunction

  // ****************************************************************************
  // FUNCTION: convert2string()
  // This function converts all variables in this class to a single string for 
  // logfile reporting.
  //
  virtual function string convert2string();
    // pragma uvmf custom convert2string begin
    // UVMF_CHANGE_ME : Customize format if desired.
    return $sformatf("read_data:0x%x write_data:0x%x address:0x%x byte_enable:0x%x chksum:0x%x ",read_data,write_data,address,byte_enable,chksum);
    // pragma uvmf custom convert2string end
  endfunction

  //*******************************************************************
  // FUNCTION: do_print()
  // This function is automatically called when the .print() function
  // is called on this class.
  //
  virtual function void do_print(uvm_printer printer);
    // pragma uvmf custom do_print begin
    // UVMF_CHANGE_ME : Current contents of do_print allows for the use of UVM 1.1d, 1.2 or P1800.2.
    // Update based on your own printing preference according to your preferred UVM version
    $display(convert2string());
    // pragma uvmf custom do_print end
  endfunction

  //*******************************************************************
  // FUNCTION: do_compare()
  // This function is automatically called when the .compare() function
  // is called on this class.
  //
  virtual function bit do_compare (uvm_object rhs, uvm_comparer comparer);
    mem_transaction #(
        .DATA_WIDTH(DATA_WIDTH),
        .ADDR_WIDTH(ADDR_WIDTH)
        ) RHS;
    if (!$cast(RHS,rhs)) return 0;
    // pragma uvmf custom do_compare begin
    // UVMF_CHANGE_ME : Eliminate comparison of variables not to be used for compare
    return (super.do_compare(rhs,comparer)
            &&(this.read_data == RHS.read_data)
            &&(this.write_data == RHS.write_data)
            &&(this.address == RHS.address)
            );
    // pragma uvmf custom do_compare end
  endfunction

  //*******************************************************************
  // FUNCTION: do_copy()
  // This function is automatically called when the .copy() function
  // is called on this class.
  //
  virtual function void do_copy (uvm_object rhs);
    mem_transaction #(
        .DATA_WIDTH(DATA_WIDTH),
        .ADDR_WIDTH(ADDR_WIDTH)
        ) RHS;
    assert($cast(RHS,rhs));
    // pragma uvmf custom do_copy begin
    super.do_copy(rhs);
    this.read_data = RHS.read_data;
    this.write_data = RHS.write_data;
    this.address = RHS.address;
    this.byte_enable = RHS.byte_enable;
    this.chksum = RHS.chksum;
    // pragma uvmf custom do_copy end
  endfunction

  // ****************************************************************************
  // FUNCTION: add_to_wave()
  // This function is used to display variables in this class in the waveform 
  // viewer.  The start_time and end_time variables must be set before this 
  // function is called.  If the start_time and end_time variables are not set
  // the transaction will be hidden at 0ns on the waveform display.
  // 
  virtual function void add_to_wave(int transaction_viewing_stream_h);
    `ifdef QUESTA
    if (transaction_view_h == 0) begin
      transaction_view_h = $begin_transaction(transaction_viewing_stream_h,"mem_transaction",start_time);
    end
    super.add_to_wave(transaction_view_h);
    // pragma uvmf custom add_to_wave begin
    // UVMF_CHANGE_ME : Color can be applied to transaction entries based on content, example below
    // case()
    //   1 : $add_color(transaction_view_h,"red");
    //   default : $add_color(transaction_view_h,"grey");
    // endcase
    // UVMF_CHANGE_ME : Eliminate transaction variables not wanted in transaction viewing in the waveform viewer
    $add_attribute(transaction_view_h,read_data,"read_data");
    $add_attribute(transaction_view_h,write_data,"write_data");
    $add_attribute(transaction_view_h,address,"address");
    $add_attribute(transaction_view_h,byte_enable,"byte_enable");
    $add_attribute(transaction_view_h,chksum,"chksum");
    // pragma uvmf custom add_to_wave end
    $end_transaction(transaction_view_h,end_time);
    $free_transaction(transaction_view_h);
    `endif // QUESTA
  endfunction

endclass

// pragma uvmf custom external begin
// pragma uvmf custom external end

